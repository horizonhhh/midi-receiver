/*
** ECE 353: Computer Systems Lab I
** Lab 4: MIDI Receiver in Verilog
**
** Ryan Lagasse, Perveshwer Jaswal, Ricardo Henriquez
*/

module HalfAdder (A, B, S, C);

endmodule

module DFlipFlop (D, CLK, Q, Qnot);

endmodule

